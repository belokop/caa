name = myPear
description = Core functions and classes for the myPear package
package = myPear
;;;
;;; Due to changes in assets treatment between different Drupal versions 
;;; this is done explicitely in myPear.module
;;;
;stylesheets[all][] = css/myPear.css
;stylesheets[all][] = css/bIcal.css
;stylesheets[all][] = css/b_table.css
;stylesheets[all][] = css/ibox.css
;stylesheets[all][] = css/drp.css

configure = admin/config/user-interface/myPear
core = 8.x
version = 3.0.3

